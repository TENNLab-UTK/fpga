`timescale 1ns/1ps

import processor_config::*;

module axis_processor_tb;

    // Simulation constants
    localparam NUM_INP = 9;

    // Simulation signals
    logic [INP_WIDTH-1:0] inp_data [0:NUM_INP-1];
    int t = 0;

    // Global signals
    logic clk;
    logic arstn;

    // AXIS master signals
    logic m_tvalid;
    logic m_tready;
    logic [OUT_WIDTH-1:0] m_tdata;
    
    // AXIS slave signals
    logic s_tvalid;
    logic s_tready;
    logic [INP_WIDTH-1:0] s_tdata;

    axis_processor uut (
        .clk(clk),
        .arstn(arstn),
        .s_axis_tdata(s_tdata),
        .s_axis_tvalid(s_tvalid),
        .s_axis_tready(s_tready),
        .m_axis_tdata(m_tdata),
        .m_axis_tvalid(m_tvalid),
        .m_axis_tready(m_tready)
    );

    // Simulate network's input data packets using AXI Stream
    initial begin: axis_inp_sim

        // inp_data[0] = 8'b10010000; // CLR, AS 0 0 1; RUN 1
        // inp_data[1] = 8'b00000100; // AS 1 0 1; RUN 1
        // inp_data[2] = 8'b00010100; // AS 0 0 1; AS 1 0 1; RUN 1
        // inp_data[3] = 8'b00000000; // RUN 1
        // inp_data[4] = 8'b00000000; // RUN 1
        // inp_data[5] = 8'b00000000; // RUN 1
        // inp_data[6] = 8'b00000000; // RUN 1
        // inp_data[7] = 8'b00000000; // RUN 1
        // inp_data[8] = 8'b01010000; // DEC; AS 0 0 1; RUN 1
        // inp_data[9] = 8'b00000100; // AS 1 0 1; RUN 1
        // inp_data[10] = 8'b00010100; // AS 0 0 1; AS 1 0 1; RUN 1
        // inp_data[11] = 8'b00000000; // RUN 1
        // inp_data[12] = 8'b00000000; // RUN 1
        // inp_data[13] = 8'b00000000; // RUN 1
        // inp_data[14] = 8'b00000000; // RUN 1
        // inp_data[15] = 8'b00000000; // RUN 1
        // inp_data[16] = 8'b01000000; // DEC; RUN 1

       inp_data[0] = 8'b01000100; // AS 0 0 1
       inp_data[1] = 8'b00100001; // RUN 1
       inp_data[2] = 8'b01010100; // AS 1 0 1
       inp_data[3] = 8'b00100001; // RUN 1
       inp_data[4] = 8'b01000100; // AS 0 0 1
       inp_data[5] = 8'b01010100; // AS 1 0 1
       inp_data[6] = 8'b00111111; // RUN 31
       inp_data[7] = 8'b00110001; // RUN 17
       inp_data[8] = 8'b10000000; // DEC
//       inp_data[10] = 8'b01000100; // AS 0 0 1
//       inp_data[11] = 8'b00100001; // RUN 1
//       inp_data[12] = 8'b01010100; // AS 1 0 1
//       inp_data[13] = 8'b00100001; // RUN 1
//       inp_data[14] = 8'b01000100; // AS 0 0 1
//       inp_data[15] = 8'b01010100; // AS 1 0 1
//       inp_data[16] = 8'b00011111; // RUN 31
//       inp_data[17] = 8'b00010001; // RUN 17
//       inp_data[18] = 8'b10000000; // DEC
        
        m_tready = 0;
        s_tvalid = 0;
        s_tdata = 0;

        // Wait for reset
        #350;

        m_tready = 1;
        #50;

        @(posedge clk);
        
        // Set valid signal high to indicate valid input packets
        s_tvalid = 1;

        // Send all input data to unit under test; for each packet, wait until a clock rising edge where s_tready is high (indicates successful AXIS handshake)
        foreach (inp_data[i]) begin
            #10;
            s_tdata = inp_data[i];
            s_tvalid = 1;
            @(posedge clk);
            while(s_tready != 1) begin
                @(posedge clk);
            end
            #10
            s_tvalid = 0;
            s_tdata = ~0;
            @(posedge clk);
        end
        
        // Set valid signal low after all input packets have been processed/sent
        #1;
        s_tvalid = 0;
    end

    // Simulate simple network's output data packet using AXI Stream
    initial begin: axis_out_sim
        forever begin
            @(posedge clk);
            if(m_tready == 1 && m_tvalid == 1) begin
                $display("%d: 0b%0b", t, m_tdata);
                t = t + 1;
            end
        end
    end

    // Simulate 10MHz clock
    initial begin: clk_sim
        clk = 0;
        forever #50 clk = ~clk;
    end

    // Simulate reset signal
    initial begin: rst_sim
        arstn = 1;
        #70;
        arstn = 0;
        #180;
        arstn = 1;
    end

endmodule: axis_processor_tb;