// Copyright (c) 2024 Keegan Dent
//
// This source describes Open Hardware and is licensed under the CERN-OHL-W v2
// You may redistribute and modify this documentation and make products using
// it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).
//
// This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED WARRANTY,
// INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY AND FITNESS FOR A
// PARTICULAR PURPOSE. Please see the CERN-OHL-W v2 for applicable conditions.

`include "macros.svh"

import processor_config::*;

module uart_processor #(
    parameter real CLK_FREQ,
    parameter int BAUD_RATE = 115_200,
    parameter int BUFFER_RX = 4096,
    parameter int BUFFER_TX = 4096
) (
    input logic clk,
    input logic arstn,
    input logic rxd,
    output logic txd,
    output logic rx_busy,
    output logic tx_busy,
    output logic rx_error
);
    // Do not change unless adding support for UART parameters outside 8N1 (likely never)
    localparam int UART_WIDTH = 8;
    localparam int UART_PADS = 2;

    logic [UART_WIDTH-1:0] rx_axis_tdata, tx_axis_tdata;
    logic rx_axis_tvalid, rx_axis_tready, tx_axis_tvalid, tx_axis_tready;
    logic rx_frame_error, rx_overrun_error;

    // This looks like odd code for a simple integer division, however
    // 1. Vivado does not seem to truncate but ROUND decimals by default, so the solution would be $floor or $rtoi
    // 2. Except Quartus won't synthesize code that uses $floor or $rtoi in even localparam math -_-
    localparam int PRESCALE = (CLK_FREQ / real'(UART_WIDTH * BAUD_RATE) - 0.5);
    logic [15:0] prescale;
    assign prescale = PRESCALE;

    uart #(
        .DATA_WIDTH(UART_WIDTH)
    ) uart_inst (
        .clk,
        .arstn,
        .s_axis_tdata(tx_axis_tdata),
        .s_axis_tvalid(tx_axis_tvalid),
        .s_axis_tready(tx_axis_tready),
        .m_axis_tdata(rx_axis_tdata),
        .m_axis_tvalid(rx_axis_tvalid),
        .m_axis_tready(rx_axis_tready),
        .rxd,
        .txd,
        .rx_busy,
        .tx_busy,
        .rx_frame_error,
        .rx_overrun_error,
        .prescale
    );

    always_ff @(posedge clk or negedge arstn) begin : set_rx_erorr
        if (arstn == 0) begin
            rx_error <= 0;
        end else begin
            rx_error <= rx_error || rx_frame_error || rx_overrun_error;
        end
    end

    logic [INP_WIDTH-1:0] inp_axis_tdata;
    logic inp_axis_tvalid, inp_axis_tready;
    logic [OUT_WIDTH-1:0] out_axis_tdata;
    logic out_axis_tvalid, out_axis_tready;

    axis_processor proc (
        .clk,
        .arstn,
        .s_axis_tdata(inp_axis_tdata),
        .s_axis_tvalid(inp_axis_tvalid),
        .s_axis_tready(inp_axis_tready),
        .m_axis_tdata(out_axis_tdata),
        .m_axis_tvalid(out_axis_tvalid),
        .m_axis_tready(out_axis_tready)
    );

    // we buffer the rx side because there is no way of conveying backpressure to the host
    // we don't buffer the tx side because the host has a buffer and the UART tx module exerts backpressure
    // the question becomes how do we size the buffer?
    // we need to anticipate how many packets we could receive while the processor is transmitting
    // - for a Dispatch Source
    //   - take the number of runs supported by the operand width (2 ^ run_width - 1)
    //   - multiply by the amount of time per run (further below)
    //   - divide by the time per packet (10 buad/byte * (out_width / 8) / baud_rate)
    // - for a Stream Source, for a Stream Source, the strategy is to mirror the size of the linux host buffer: 4096 bytes
    // the worst case run latency is driven by the UART baud rate, the system clock speed, and the sink mechanism
    // for Dispatch Sink it's the sum of:
    // - one clock per net_out
    // - ten baud per byte; max_bytes is (net_out + 1) * (out_width / 8)
    // for Stream Sink it's again ten baud per byte; max_bytes is (out_width / 8)
    // clock cycle per bit actually transmitted, rounded up
    localparam int CLK_PER_BIT = CLK_FREQ / (UART_WIDTH * BAUD_RATE / (UART_WIDTH + UART_PADS)) + 0.5;
    // number of
    localparam int BIT_PER_RUN_MAX = OUT_PER_RUN_MAX * OUT_WIDTH;
    localparam int CLK_PER_RUN_MAX = CLK_PER_BIT * BIT_PER_RUN_MAX + OUT_PER_RUN_MAX - 1;
    localparam int RUN_MAX = `min(RUN_MAX_BASE ** RUN_WIDTH - 1, `width_bytes_to_bits(BUFFER_RX) / BIT_PER_RUN_MAX);
    localparam int CLK_MAX = CLK_PER_RUN_MAX * RUN_MAX;
    localparam int BUF_BYTES = `max(BUFFER_RX, `width_bits_to_bytes(CLK_MAX / CLK_PER_BIT));

    logic [UART_WIDTH-1:0] buf_axis_tdata;
    logic buf_axis_tvalid, buf_axis_tready;

    axis_pipeline_register #(
        .DATA_WIDTH(UART_WIDTH),
        .LENGTH(BUF_BYTES)
    ) rx_buf (
        .clk,
        .arstn,
        .s_axis_tdata(rx_axis_tdata),
        .s_axis_tvalid(rx_axis_tvalid),
        .s_axis_tready(rx_axis_tready),
        .m_axis_tdata(buf_axis_tdata),
        .m_axis_tvalid(buf_axis_tvalid),
        .m_axis_tready(buf_axis_tready)
    );

    axis_adapter #(
        .S_DATA_WIDTH(UART_WIDTH),
        .S_KEEP_ENABLE(0),
        .M_DATA_WIDTH(INP_WIDTH),
        .M_KEEP_ENABLE(0)
    )  rx_inp_adapter (
        .clk,
        .arstn,
        .s_axis_tdata(buf_axis_tdata),
        .s_axis_tvalid(buf_axis_tvalid),
        .s_axis_tready(buf_axis_tready),
        .m_axis_tdata(inp_axis_tdata),
        .m_axis_tvalid(inp_axis_tvalid),
        .m_axis_tready(inp_axis_tready)
    );

    axis_adapter #(
        .S_DATA_WIDTH(OUT_WIDTH),
        .S_KEEP_ENABLE(0),
        .M_DATA_WIDTH(UART_WIDTH),
        .M_KEEP_ENABLE(0)
    ) out_tx_adapter (
        .clk,
        .arstn,
        .s_axis_tdata(out_axis_tdata),
        .s_axis_tvalid(out_axis_tvalid),
        .s_axis_tready(out_axis_tready),
        .m_axis_tdata(tx_axis_tdata),
        .m_axis_tvalid(tx_axis_tvalid),
        .m_axis_tready(tx_axis_tready)
    );
endmodule
