`timescale 1ns/1ps

import processor_tlast_config::*;

module dma_simple_axis_tb;

    // Simulation constants
    localparam NUM_INP = 131;

    // Simulation signals
    logic [(INP_TDATA_WIDTH_BYTES * 8 - 1):0] inp_data [0:NUM_INP-1];
    int t = 0;

    // Global signals
    logic clk;
    logic arstn;

    // AXIS master signals
    logic m_tvalid;
    logic m_tready;
    logic [(OUT_TDATA_WIDTH_BYTES * 8 - 1):0] m_tdata;
    logic [OUT_TDATA_WIDTH_BYTES-1:0] m_tkeep;
    logic m_tlast;
    
    // AXIS slave signals
    logic s_tvalid;
    logic s_tready;
    logic [(INP_TDATA_WIDTH_BYTES * 8 - 1):0] s_tdata;
    logic [INP_TDATA_WIDTH_BYTES-1:0] s_tkeep;
    logic s_tlast;

    axis #(.DATA_WIDTH_BYTES(INP_TDATA_WIDTH_BYTES)) s_axis();
    axis #(.DATA_WIDTH_BYTES(OUT_TDATA_WIDTH_BYTES)) m_axis();

    assign s_axis.tvalid = s_tvalid;
    assign s_tready = s_axis.tready;
    assign s_axis.tdata = s_tdata;
    assign s_axis.tkeep = s_tkeep;
    assign s_axis.tlast = s_tlast;
    assign m_tvalid = m_axis.tvalid;
    assign m_axis.tready = m_tready;
    assign m_tdata = m_axis.tdata;
    assign m_tkeep = m_axis.tkeep;
    assign m_tlast = m_axis.tlast;

    axis_processor_tlast uut (
        .clk(clk),
        .arstn(arstn),
        .s_axis(s_axis),
        .m_axis(m_axis)
    );

    // Simulate simple network's input data packet using AXI Stream
    initial begin: axis_inp_sim


        // Fill test input array with input pkts
        inp_data[0] = 64'b0000000000000000000000000000000000010000100000000000000000000000;
        inp_data[1] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[2] = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        inp_data[3] = 64'b0000000000000000000000000100000000000000000001000000000000000000;
        inp_data[4] = 64'b0000000000000001000000000000000000000000000000000000000000000000;
        inp_data[5] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[6] = 64'b0000010000100000000000000000000000000000000000000000000000000000;
        inp_data[7] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[8] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[9] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[10] = 64'b0000000000100000000000000000000000000000000000000000000000000000;
        inp_data[11] = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        inp_data[12] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[13] = 64'b0000000000000000000000000000000000010000000001000000000000000000;
        inp_data[14] = 64'b0000000000000001000000000000000000000000000001000000000000000000;
        inp_data[15] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[16] = 64'b0000010000100000000000000000000000000000000000000000000000000000;
        inp_data[17] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[18] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[19] = 64'b0000000000000001000000000000000000000000100000000000000000000000;
        inp_data[20] = 64'b0000010000000000000000000100000000000000000000000000000000000000;
        inp_data[21] = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        inp_data[22] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[23] = 64'b0000000000000000000010000000000000000000000001000000000000000000;
        inp_data[24] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[25] = 64'b0000000000000000000010000100000000000000000000000000000000000000;
        inp_data[26] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[27] = 64'b0000000000000001000000000000000000000000000000000000000000000000;
        inp_data[28] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[29] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[30] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[31] = 64'b0000000000000000000000000100000000000000000001000000000000000000;
        inp_data[32] = 64'b0000000000100000000000000000001000010000000000000000000000000000;
        inp_data[33] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[34] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[35] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[36] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[37] = 64'b0000000000000000000010000000000000000000000000000000000000000000;
        inp_data[38] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[39] = 64'b0000000000000000000000000000000000000000100000000000000000000000;
        inp_data[40] = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        inp_data[41] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[42] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[43] = 64'b0000000000000001000000000000000000000000000000000000000000000000;
        inp_data[44] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[45] = 64'b0000000000000000000000000000001000000000000001000000000000000000;
        inp_data[46] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[47] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[48] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[49] = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        inp_data[50] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[51] = 64'b0000010000000001000000000000001000000000100000000000000000000000;
        inp_data[52] = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        inp_data[53] = 64'b0000000000000000000000000100000000000000000000000000000000000000;
        inp_data[54] = 64'b0000000000000000000000000000000000000000100000000000000000000000;
        inp_data[55] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[56] = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        inp_data[57] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[58] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[59] = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        inp_data[60] = 64'b0000000000000001000000000000000000000000000000000000000000000000;
        inp_data[61] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[62] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[63] = 64'b0000000000000000000010000000000000000000000000000000000000000000;
        inp_data[64] = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        inp_data[65] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[66] = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        inp_data[67] = 64'b0000000000100000000000000000000000000000000000000000000000000000;
        inp_data[68] = 64'b0000000000000001000000000000000000000000000000000000000000000000;
        inp_data[69] = 64'b0000000000000001000000000000001000000000000000000000000000000000;
        inp_data[70] = 64'b0000010000000000000000000000000000000000000001000000000000000000;
        inp_data[71] = 64'b0000000000000000000010000000000000000000000000000000000000000000;
        inp_data[72] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[73] = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        inp_data[74] = 64'b0000010000000001000010000000000000000000000000000000000000000000;
        inp_data[75] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[76] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[77] = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        inp_data[78] = 64'b0000000000000001000000000000000000000000100000000000000000000000;
        inp_data[79] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[80] = 64'b0000000000000000000000000100000000000000000000000000000000000000;
        inp_data[81] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[82] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[83] = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        inp_data[84] = 64'b0000000000000001000000000000000000000000100000000000000000000000;
        inp_data[85] = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        inp_data[86] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[87] = 64'b0000000000000000000000000000000000000000100000000000000000000000;
        inp_data[88] = 64'b0000000000000000000000000000000000000000100000000000000000000000;
        inp_data[89] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[90] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[91] = 64'b0000000000000000000000000100000000000000000000000000000000000000;
        inp_data[92] = 64'b0000010000000000000000000000000000000000100000000000000000000000;
        inp_data[93] = 64'b0000000000000000000010000000000000000000100000000000000000000000;
        inp_data[94] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[95] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[96] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[97] = 64'b0000000000000000000000000100000000000000000000000000000000000000;
        inp_data[98] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[99] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[100] = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        inp_data[101] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[102] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[103] = 64'b0000010000000000000000000000000000000000100000000000000000000000;
        inp_data[104] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[105] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[106] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[107] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[108] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[109] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[110] = 64'b0000000000100000000010000000000000010000000000000000000000000000;
        inp_data[111] = 64'b0000010000100000000010000100000000000000000000000000000000000000;
        inp_data[112] = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        inp_data[113] = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        inp_data[114] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[115] = 64'b0000000000100000000010000000000000000000000000000000000000000000;
        inp_data[116] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[117] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[118] = 64'b0000010000000000000000000000001000010000000000000000000000000000;
        inp_data[119] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[120] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[121] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[122] = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        inp_data[123] = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        inp_data[124] = 64'b0000000000100000000000000000001000000000100000000000000000000000;
        inp_data[125] = 64'b0000000000000000000010000000000000000000100000000000000000000000;
        inp_data[126] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[127] = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        inp_data[128] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[129] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        inp_data[130] = 64'b0000000000000000000000000000000000000000000000000000000000000000;


        
        m_tready = 0;
        s_tvalid = 0;
        s_tdata = 0;
        s_tkeep = 0;
        s_tlast = 0;

        // Wait for reset
        #350;

        // Assign m_tready to high for the whole simulation
        m_tready = 1;
        #50;

        @(posedge clk);

        // Set valid input data packet and 
        
        // Set valid and all tkeep signals high to indicate valid input packets
        s_tkeep = ~0;
        s_tvalid = 1;

        // Send all input data to unit under test; for each packet, wait until a clock rising edge where s_tready is high (indicates successful AXIS handshake)
        foreach (inp_data[i]) begin
            s_tdata = inp_data[i];
            @(posedge clk);
            while(s_tready != 1) begin
                @(posedge clk);
            end
        end
        
        s_tvalid = 0;
    end

    // Simulate simple network's output data packet using AXI Stream
    initial begin: axis_out_sim
        forever begin
            @(posedge clk);
            if(m_tready == 1 && m_tvalid == 1) begin
                $display("%d: 0b%0b", t, m_tdata);
                t = t + 1;
            end
        end
    end

    // Simulate 10MHz clock
    initial begin: clk_sim
        clk = 0;
        forever #50 clk = ~clk;
    end

    // Simulate reset signal
    initial begin: rst_sim
        arstn = 1;
        #70;
        arstn = 0;
        #180;
        arstn = 1;
    end

endmodule: dma_simple_axis_tb;